magic
tech sky130A
magscale 1 2
timestamp 1764449767
<< pwell >>
rect -404 -728 404 728
<< nmos >>
rect -208 318 -108 518
rect -50 318 50 518
rect 108 318 208 518
rect -208 -100 -108 100
rect -50 -100 50 100
rect 108 -100 208 100
rect -208 -518 -108 -318
rect -50 -518 50 -318
rect 108 -518 208 -318
<< ndiff >>
rect -266 506 -208 518
rect -266 330 -254 506
rect -220 330 -208 506
rect -266 318 -208 330
rect -108 506 -50 518
rect -108 330 -96 506
rect -62 330 -50 506
rect -108 318 -50 330
rect 50 506 108 518
rect 50 330 62 506
rect 96 330 108 506
rect 50 318 108 330
rect 208 506 266 518
rect 208 330 220 506
rect 254 330 266 506
rect 208 318 266 330
rect -266 88 -208 100
rect -266 -88 -254 88
rect -220 -88 -208 88
rect -266 -100 -208 -88
rect -108 88 -50 100
rect -108 -88 -96 88
rect -62 -88 -50 88
rect -108 -100 -50 -88
rect 50 88 108 100
rect 50 -88 62 88
rect 96 -88 108 88
rect 50 -100 108 -88
rect 208 88 266 100
rect 208 -88 220 88
rect 254 -88 266 88
rect 208 -100 266 -88
rect -266 -330 -208 -318
rect -266 -506 -254 -330
rect -220 -506 -208 -330
rect -266 -518 -208 -506
rect -108 -330 -50 -318
rect -108 -506 -96 -330
rect -62 -506 -50 -330
rect -108 -518 -50 -506
rect 50 -330 108 -318
rect 50 -506 62 -330
rect 96 -506 108 -330
rect 50 -518 108 -506
rect 208 -330 266 -318
rect 208 -506 220 -330
rect 254 -506 266 -330
rect 208 -518 266 -506
<< ndiffc >>
rect -254 330 -220 506
rect -96 330 -62 506
rect 62 330 96 506
rect 220 330 254 506
rect -254 -88 -220 88
rect -96 -88 -62 88
rect 62 -88 96 88
rect 220 -88 254 88
rect -254 -506 -220 -330
rect -96 -506 -62 -330
rect 62 -506 96 -330
rect 220 -506 254 -330
<< psubdiff >>
rect -368 658 -272 692
rect 272 658 368 692
rect -368 596 -334 658
rect 334 596 368 658
rect -368 -658 -334 -596
rect 334 -658 368 -596
rect -368 -692 -272 -658
rect 272 -692 368 -658
<< psubdiffcont >>
rect -272 658 272 692
rect -368 -596 -334 596
rect 334 -596 368 596
rect -272 -692 272 -658
<< poly >>
rect -208 590 -108 606
rect -208 556 -192 590
rect -124 556 -108 590
rect -208 518 -108 556
rect -50 590 50 606
rect -50 556 -34 590
rect 34 556 50 590
rect -50 518 50 556
rect 108 590 208 606
rect 108 556 124 590
rect 192 556 208 590
rect 108 518 208 556
rect -208 280 -108 318
rect -208 246 -192 280
rect -124 246 -108 280
rect -208 230 -108 246
rect -50 280 50 318
rect -50 246 -34 280
rect 34 246 50 280
rect -50 230 50 246
rect 108 280 208 318
rect 108 246 124 280
rect 192 246 208 280
rect 108 230 208 246
rect -208 172 -108 188
rect -208 138 -192 172
rect -124 138 -108 172
rect -208 100 -108 138
rect -50 172 50 188
rect -50 138 -34 172
rect 34 138 50 172
rect -50 100 50 138
rect 108 172 208 188
rect 108 138 124 172
rect 192 138 208 172
rect 108 100 208 138
rect -208 -138 -108 -100
rect -208 -172 -192 -138
rect -124 -172 -108 -138
rect -208 -188 -108 -172
rect -50 -138 50 -100
rect -50 -172 -34 -138
rect 34 -172 50 -138
rect -50 -188 50 -172
rect 108 -138 208 -100
rect 108 -172 124 -138
rect 192 -172 208 -138
rect 108 -188 208 -172
rect -208 -246 -108 -230
rect -208 -280 -192 -246
rect -124 -280 -108 -246
rect -208 -318 -108 -280
rect -50 -246 50 -230
rect -50 -280 -34 -246
rect 34 -280 50 -246
rect -50 -318 50 -280
rect 108 -246 208 -230
rect 108 -280 124 -246
rect 192 -280 208 -246
rect 108 -318 208 -280
rect -208 -556 -108 -518
rect -208 -590 -192 -556
rect -124 -590 -108 -556
rect -208 -606 -108 -590
rect -50 -556 50 -518
rect -50 -590 -34 -556
rect 34 -590 50 -556
rect -50 -606 50 -590
rect 108 -556 208 -518
rect 108 -590 124 -556
rect 192 -590 208 -556
rect 108 -606 208 -590
<< polycont >>
rect -192 556 -124 590
rect -34 556 34 590
rect 124 556 192 590
rect -192 246 -124 280
rect -34 246 34 280
rect 124 246 192 280
rect -192 138 -124 172
rect -34 138 34 172
rect 124 138 192 172
rect -192 -172 -124 -138
rect -34 -172 34 -138
rect 124 -172 192 -138
rect -192 -280 -124 -246
rect -34 -280 34 -246
rect 124 -280 192 -246
rect -192 -590 -124 -556
rect -34 -590 34 -556
rect 124 -590 192 -556
<< locali >>
rect -368 658 -272 692
rect 272 658 368 692
rect -368 596 -334 658
rect 334 596 368 658
rect -237 556 -192 590
rect -124 556 -34 590
rect 34 556 124 590
rect 192 556 237 590
rect -254 506 -220 522
rect -254 314 -220 330
rect -96 506 -62 522
rect -96 314 -62 330
rect 62 506 96 522
rect 62 314 96 330
rect 220 506 254 522
rect 220 314 254 330
rect -237 246 -192 280
rect -124 246 -34 280
rect 34 246 124 280
rect 192 246 237 280
rect -237 138 -192 172
rect -124 138 -34 172
rect 34 138 124 172
rect 192 138 237 172
rect -254 88 -220 104
rect -254 -104 -220 -88
rect -96 88 -62 104
rect -96 -104 -62 -88
rect 62 88 96 104
rect 62 -104 96 -88
rect 220 88 254 104
rect 220 -104 254 -88
rect -237 -172 -192 -138
rect -124 -172 -34 -138
rect 34 -172 124 -138
rect 192 -172 237 -138
rect -237 -280 -192 -246
rect -124 -280 -34 -246
rect 34 -280 124 -246
rect 192 -280 237 -246
rect -254 -330 -220 -314
rect -254 -522 -220 -506
rect -96 -330 -62 -314
rect -96 -522 -62 -506
rect 62 -330 96 -314
rect 62 -522 96 -506
rect 220 -330 254 -314
rect 220 -522 254 -506
rect -237 -590 -192 -556
rect -124 -590 -34 -556
rect 34 -590 124 -556
rect 192 -590 237 -556
rect -368 -658 -334 -596
rect 334 -658 368 -596
rect -368 -692 -272 -658
rect 272 -692 368 -658
<< viali >>
rect -192 556 -124 590
rect -34 556 34 590
rect 124 556 192 590
rect -254 330 -220 506
rect -96 330 -62 506
rect 62 330 96 506
rect 220 330 254 506
rect -192 246 -124 280
rect -34 246 34 280
rect 124 246 192 280
rect -192 138 -124 172
rect -34 138 34 172
rect 124 138 192 172
rect -254 -88 -220 88
rect -96 -88 -62 88
rect 62 -88 96 88
rect 220 -88 254 88
rect -192 -172 -124 -138
rect -34 -172 34 -138
rect 124 -172 192 -138
rect -192 -280 -124 -246
rect -34 -280 34 -246
rect 124 -280 192 -246
rect -254 -506 -220 -330
rect -96 -506 -62 -330
rect 62 -506 96 -330
rect 220 -506 254 -330
rect -192 -590 -124 -556
rect -34 -590 34 -556
rect 124 -590 192 -556
<< metal1 >>
rect -204 590 -112 596
rect -46 590 46 596
rect 112 590 204 596
rect -237 556 -192 590
rect -124 556 -34 590
rect 34 556 124 590
rect 192 556 237 590
rect -204 550 -112 556
rect -46 550 46 556
rect 112 550 204 556
rect -260 506 -214 518
rect -260 330 -254 506
rect -220 330 -214 506
rect -260 318 -214 330
rect -102 506 -56 518
rect -102 330 -96 506
rect -62 330 -56 506
rect -102 318 -56 330
rect 56 506 102 518
rect 56 330 62 506
rect 96 330 102 506
rect 56 318 102 330
rect 214 506 260 518
rect 214 330 220 506
rect 254 330 260 506
rect 214 318 260 330
rect -204 280 -112 286
rect -46 280 46 286
rect 112 280 204 286
rect -237 246 -192 280
rect -124 246 -34 280
rect 34 246 124 280
rect 192 246 237 280
rect -204 240 -112 246
rect -46 240 46 246
rect 112 240 204 246
rect -204 172 -112 178
rect -46 172 46 178
rect 112 172 204 178
rect -237 138 -192 172
rect -124 138 -34 172
rect 34 138 124 172
rect 192 138 237 172
rect -204 132 -112 138
rect -46 132 46 138
rect 112 132 204 138
rect -260 88 -214 100
rect -260 -88 -254 88
rect -220 -88 -214 88
rect -260 -100 -214 -88
rect -102 88 -56 100
rect -102 -88 -96 88
rect -62 -88 -56 88
rect -102 -100 -56 -88
rect 56 88 102 100
rect 56 -88 62 88
rect 96 -88 102 88
rect 56 -100 102 -88
rect 214 88 260 100
rect 214 -88 220 88
rect 254 -88 260 88
rect 214 -100 260 -88
rect -204 -138 -112 -132
rect -46 -138 46 -132
rect 112 -138 204 -132
rect -237 -172 -192 -138
rect -124 -172 -34 -138
rect 34 -172 124 -138
rect 192 -172 237 -138
rect -204 -178 -112 -172
rect -46 -178 46 -172
rect 112 -178 204 -172
rect -204 -246 -112 -240
rect -46 -246 46 -240
rect 112 -246 204 -240
rect -237 -280 -192 -246
rect -124 -280 -34 -246
rect 34 -280 124 -246
rect 192 -280 237 -246
rect -204 -286 -112 -280
rect -46 -286 46 -280
rect 112 -286 204 -280
rect -260 -330 -214 -318
rect -260 -506 -254 -330
rect -220 -506 -214 -330
rect -260 -518 -214 -506
rect -102 -330 -56 -318
rect -102 -506 -96 -330
rect -62 -506 -56 -330
rect -102 -518 -56 -506
rect 56 -330 102 -318
rect 56 -506 62 -330
rect 96 -506 102 -330
rect 56 -518 102 -506
rect 214 -330 260 -318
rect 214 -506 220 -330
rect 254 -506 260 -330
rect 214 -518 260 -506
rect -204 -556 -112 -550
rect -46 -556 46 -550
rect 112 -556 204 -550
rect -237 -590 -192 -556
rect -124 -590 -34 -556
rect 34 -590 124 -556
rect 192 -590 237 -556
rect -204 -596 -112 -590
rect -46 -596 46 -590
rect 112 -596 204 -590
<< labels >>
rlabel psubdiffcont 0 -675 0 -675 0 B
port 17 nsew
rlabel ndiffc -237 -418 -237 -418 0 D0_0
port 18 nsew
rlabel polycont -158 -263 -158 -263 0 G0
port 3 nsew
rlabel ndiffc -237 0 -237 0 0 D0_1
port 19 nsew
rlabel polycont -158 155 -158 155 0 G1
port 5 nsew
rlabel ndiffc -237 418 -237 418 0 D0_2
port 20 nsew
rlabel polycont -158 573 -158 573 0 G2
port 7 nsew
rlabel ndiffc -79 -418 -79 -418 0 S1_0
port 21 nsew
rlabel polycont 0 -263 0 -263 0 G0
port 3 nsew
rlabel ndiffc -79 0 -79 0 0 S1_1
port 22 nsew
rlabel polycont 0 155 0 155 0 G1
port 5 nsew
rlabel ndiffc -79 418 -79 418 0 S1_2
port 23 nsew
rlabel polycont 0 573 0 573 0 G2
port 7 nsew
rlabel ndiffc 79 -418 79 -418 0 D2_0
port 24 nsew
rlabel ndiffc 237 -418 237 -418 0 S2_0
port 25 nsew
rlabel polycont 158 -263 158 -263 0 G0
port 3 nsew
rlabel ndiffc 79 0 79 0 0 D2_1
port 26 nsew
rlabel ndiffc 237 0 237 0 0 S2_1
port 27 nsew
rlabel polycont 158 155 158 155 0 G1
port 5 nsew
rlabel ndiffc 79 418 79 418 0 D2_2
port 28 nsew
rlabel ndiffc 237 418 237 418 0 S2_2
port 29 nsew
rlabel polycont 158 573 158 573 0 G2
port 7 nsew
<< properties >>
string FIXED_BBOX -351 -675 351 675
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.5 m 3 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
