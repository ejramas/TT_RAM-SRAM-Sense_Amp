magic
tech sky130A
magscale 1 2
timestamp 1764192597
<< error_p >>
rect -29 9281 29 9287
rect -29 9247 -17 9281
rect -29 9241 29 9247
rect -29 -9247 29 -9241
rect -29 -9281 -17 -9247
rect -29 -9287 29 -9281
<< nwell >>
rect -214 -9419 214 9419
<< pmos >>
rect -18 -9200 18 9200
<< pdiff >>
rect -76 9188 -18 9200
rect -76 -9188 -64 9188
rect -30 -9188 -18 9188
rect -76 -9200 -18 -9188
rect 18 9188 76 9200
rect 18 -9188 30 9188
rect 64 -9188 76 9188
rect 18 -9200 76 -9188
<< pdiffc >>
rect -64 -9188 -30 9188
rect 30 -9188 64 9188
<< nsubdiff >>
rect -178 9349 -82 9383
rect 82 9349 178 9383
rect -178 9287 -144 9349
rect 144 9287 178 9349
rect -178 -9349 -144 -9287
rect 144 -9349 178 -9287
rect -178 -9383 -82 -9349
rect 82 -9383 178 -9349
<< nsubdiffcont >>
rect -82 9349 82 9383
rect -178 -9287 -144 9287
rect 144 -9287 178 9287
rect -82 -9383 82 -9349
<< poly >>
rect -33 9281 33 9297
rect -33 9247 -17 9281
rect 17 9247 33 9281
rect -33 9231 33 9247
rect -18 9200 18 9231
rect -18 -9231 18 -9200
rect -33 -9247 33 -9231
rect -33 -9281 -17 -9247
rect 17 -9281 33 -9247
rect -33 -9297 33 -9281
<< polycont >>
rect -17 9247 17 9281
rect -17 -9281 17 -9247
<< locali >>
rect -178 9349 -82 9383
rect 82 9349 178 9383
rect -178 9287 -144 9349
rect 144 9287 178 9349
rect -33 9247 -17 9281
rect 17 9247 33 9281
rect -64 9188 -30 9204
rect -64 -9204 -30 -9188
rect 30 9188 64 9204
rect 30 -9204 64 -9188
rect -33 -9281 -17 -9247
rect 17 -9281 33 -9247
rect -178 -9349 -144 -9287
rect 144 -9349 178 -9287
rect -178 -9383 -82 -9349
rect 82 -9383 178 -9349
<< viali >>
rect -17 9247 17 9281
rect -64 -9188 -30 9188
rect 30 -9188 64 9188
rect -17 -9281 17 -9247
<< metal1 >>
rect -29 9281 29 9287
rect -29 9247 -17 9281
rect 17 9247 29 9281
rect -29 9241 29 9247
rect -70 9188 -24 9200
rect -70 -9188 -64 9188
rect -30 -9188 -24 9188
rect -70 -9200 -24 -9188
rect 24 9188 70 9200
rect 24 -9188 30 9188
rect 64 -9188 70 9188
rect 24 -9200 70 -9188
rect -29 -9247 29 -9241
rect -29 -9281 -17 -9247
rect 17 -9281 29 -9247
rect -29 -9287 29 -9281
<< labels >>
rlabel nsubdiffcont 0 -9366 0 -9366 0 B
port 5 nsew
rlabel pdiffc -47 0 -47 0 0 D
port 6 nsew
rlabel pdiffc 47 0 47 0 0 S
port 7 nsew
rlabel polycont 0 9264 0 9264 0 G
port 8 nsew
<< properties >>
string FIXED_BBOX -161 -9366 161 9366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 92 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
