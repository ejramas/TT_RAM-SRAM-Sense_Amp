magic
tech sky130A
magscale 1 2
timestamp 1764206135
<< error_p >>
rect 3102 11772 3108 11778
rect 3012 11771 3114 11772
rect 3107 11766 3114 11771
rect 3107 11546 3108 11766
rect 3107 11541 3114 11546
rect 3012 11540 3114 11541
rect 3102 11534 3108 11540
<< error_s >>
rect 1006 18770 1086 18778
rect 132 18647 190 18653
rect 132 18613 144 18647
rect 843 18640 901 18646
rect 132 18607 190 18613
rect 843 18606 855 18640
rect 843 18600 901 18606
rect -654 17126 -652 17196
rect 1260 13660 1340 18770
rect 1428 17151 1450 18551
rect 1456 17123 1478 18579
rect 1534 17123 1560 18579
rect 1562 17151 1588 18551
rect 1428 15515 1450 16915
rect 1456 15487 1478 16943
rect 1534 15487 1560 16943
rect 1562 15515 1588 16915
rect 1428 13879 1450 15279
rect 1456 13851 1478 15307
rect 1534 13851 1560 15307
rect 1562 13879 1588 15279
rect 1428 13026 1450 13426
rect 1456 12998 1478 13454
rect 1534 12998 1560 13454
rect 1562 13026 1588 13426
rect 1428 12408 1450 12808
rect 1456 12380 1478 12836
rect 1534 12380 1560 12836
rect 1562 12408 1588 12808
rect 1428 11790 1450 12190
rect 1456 11762 1478 12218
rect 1534 11762 1560 12218
rect 1562 11790 1588 12190
rect 2818 11772 2824 11778
rect 2812 11771 3012 11772
rect 2812 11766 2819 11771
rect 2818 11546 2819 11766
rect 2812 11541 2819 11546
rect 2812 11540 3012 11541
rect 2818 11534 2824 11540
rect 1430 6526 1450 6926
rect 1458 6498 1478 6954
rect 1534 6498 1560 6954
rect 1562 6526 1588 6926
rect 1430 5908 1450 6308
rect 1458 5880 1478 6336
rect 1534 5880 1560 6336
rect 1562 5908 1588 6308
rect 1006 5050 1086 5304
rect 1430 5290 1450 5690
rect 1458 5262 1478 5718
rect 1534 5262 1560 5718
rect 1562 5290 1588 5690
rect 91 166 137 172
rect 185 166 231 172
rect 802 159 848 172
rect 896 159 942 172
rect 116 138 259 144
rect 774 131 930 144
rect 1260 -60 1340 5050
rect 1430 3431 1450 4831
rect 1458 3403 1478 4859
rect 1534 3403 1560 4859
rect 1562 3431 1588 4831
rect 1430 1795 1450 3195
rect 1458 1767 1478 3223
rect 1534 1767 1560 3223
rect 1562 1795 1588 3195
rect 1430 159 1450 1559
rect 1458 131 1478 1587
rect 1534 131 1560 1587
rect 1562 159 1588 1559
<< metal1 >>
rect 1456 11690 1560 18998
rect 1840 7140 1900 18980
rect 1458 7040 1900 7140
rect 116 54 930 144
rect 1458 58 1560 7040
<< metal2 >>
rect 1560 11790 1620 18580
rect 1552 11702 1620 11790
rect 1560 11440 1620 11702
rect 1460 11380 1620 11440
rect 1460 10860 1560 11380
rect 1560 140 1620 6940
<< metal3 >>
rect 1400 10860 1460 13420
<< via3 >>
rect 2818 11540 3108 11772
use sky130_fd_pr__nfet_01v8_5Y7G3K  sky130_fd_pr__nfet_01v8_5Y7G3K_0
timestamp 1764192597
transform 1 0 1506 0 1 7570
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_KXEGWR  sky130_fd_pr__nfet_01v8_KXEGWR_0
timestamp 1764206135
transform 1 0 1500 0 1 11081
box -187 -288 187 288
use sky130_fd_pr__nfet_01v8_VGHGWH  sky130_fd_pr__nfet_01v8_VGHGWH_0
timestamp 1764195345
transform 1 0 1506 0 1 12608
box -246 -1028 246 1028
use sky130_fd_pr__nfet_01v8_VGHGWH  sky130_fd_pr__nfet_01v8_VGHGWH_1
timestamp 1764195345
transform 1 0 1506 0 1 6108
box -246 -1028 246 1028
use sky130_fd_pr__pfet_01v8_KT2VVS  sky130_fd_pr__pfet_01v8_KT2VVS_0
timestamp 1764192597
transform 1 0 161 0 1 9366
box -214 -9419 214 9419
use sky130_fd_pr__pfet_01v8_KT2VVS  sky130_fd_pr__pfet_01v8_KT2VVS_1
timestamp 1764192597
transform 1 0 872 0 1 9359
box -214 -9419 214 9419
use sky130_fd_pr__pfet_01v8_QGVNTY  sky130_fd_pr__pfet_01v8_QGVNTY_0
timestamp 1764202196
transform 1 0 1506 0 -1 16215
box -246 -2555 246 2555
use sky130_fd_pr__pfet_01v8_QGVNTY  sky130_fd_pr__pfet_01v8_QGVNTY_1
timestamp 1764202196
transform 1 0 1506 0 -1 2495
box -246 -2555 246 2555
use sky130_fd_pr__res_xhigh_po_0p35_RZH895  sky130_fd_pr__res_xhigh_po_0p35_RZH895_0
timestamp 1764189913
transform 0 1 -688 -1 0 17161
box -201 -632 201 632
<< end >>
