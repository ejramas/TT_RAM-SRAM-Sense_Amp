magic
tech sky130A
magscale 1 2
timestamp 1764192597
<< pwell >>
rect -246 -410 246 410
<< nmos >>
rect -50 -200 50 200
<< ndiff >>
rect -108 188 -50 200
rect -108 -188 -96 188
rect -62 -188 -50 188
rect -108 -200 -50 -188
rect 50 188 108 200
rect 50 -188 62 188
rect 96 -188 108 188
rect 50 -200 108 -188
<< ndiffc >>
rect -96 -188 -62 188
rect 62 -188 96 188
<< psubdiff >>
rect -210 340 -114 374
rect 114 340 210 374
rect -210 278 -176 340
rect 176 278 210 340
rect -210 -340 -176 -278
rect 176 -340 210 -278
rect -210 -374 -114 -340
rect 114 -374 210 -340
<< psubdiffcont >>
rect -114 340 114 374
rect -210 -278 -176 278
rect 176 -278 210 278
rect -114 -374 114 -340
<< poly >>
rect -50 272 50 288
rect -50 238 -34 272
rect 34 238 50 272
rect -50 200 50 238
rect -50 -238 50 -200
rect -50 -272 -34 -238
rect 34 -272 50 -238
rect -50 -288 50 -272
<< polycont >>
rect -34 238 34 272
rect -34 -272 34 -238
<< locali >>
rect -210 340 -114 374
rect 114 340 210 374
rect -210 278 -176 340
rect 176 278 210 340
rect -50 238 -34 272
rect 34 238 50 272
rect -96 188 -62 204
rect -96 -204 -62 -188
rect 62 188 96 204
rect 62 -204 96 -188
rect -50 -272 -34 -238
rect 34 -272 50 -238
rect -210 -340 -176 -278
rect 176 -340 210 -278
rect -210 -374 -114 -340
rect 114 -374 210 -340
<< viali >>
rect -34 238 34 272
rect -96 -188 -62 188
rect 62 -188 96 188
rect -34 -272 34 -238
<< metal1 >>
rect -46 272 46 278
rect -46 238 -34 272
rect 34 238 46 272
rect -46 232 46 238
rect -102 188 -56 200
rect -102 -188 -96 188
rect -62 -188 -56 188
rect -102 -200 -56 -188
rect 56 188 102 200
rect 56 -188 62 188
rect 96 -188 102 188
rect 56 -200 102 -188
rect -46 -238 46 -232
rect -46 -272 -34 -238
rect 34 -272 46 -238
rect -46 -278 46 -272
<< labels >>
rlabel psubdiffcont 0 -357 0 -357 0 B
port 13 nsew
rlabel ndiffc -79 0 -79 0 0 D
port 14 nsew
rlabel ndiffc 79 0 79 0 0 S
port 15 nsew
rlabel polycont 0 255 0 255 0 G
port 16 nsew
<< properties >>
string FIXED_BBOX -193 -357 193 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
