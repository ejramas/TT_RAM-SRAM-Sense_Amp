magic
tech sky130A
magscale 1 2
timestamp 1764449767
<< nwell >>
rect -214 -1219 214 1219
<< pmos >>
rect -18 -1000 18 1000
<< pdiff >>
rect -76 988 -18 1000
rect -76 -988 -64 988
rect -30 -988 -18 988
rect -76 -1000 -18 -988
rect 18 988 76 1000
rect 18 -988 30 988
rect 64 -988 76 988
rect 18 -1000 76 -988
<< pdiffc >>
rect -64 -988 -30 988
rect 30 -988 64 988
<< nsubdiff >>
rect -178 1149 -82 1183
rect 82 1149 178 1183
rect -178 1087 -144 1149
rect 144 1087 178 1149
rect -178 -1149 -144 -1087
rect 144 -1149 178 -1087
rect -178 -1183 -82 -1149
rect 82 -1183 178 -1149
<< nsubdiffcont >>
rect -82 1149 82 1183
rect -178 -1087 -144 1087
rect 144 -1087 178 1087
rect -82 -1183 82 -1149
<< poly >>
rect -33 1081 33 1097
rect -33 1047 -17 1081
rect 17 1047 33 1081
rect -33 1031 33 1047
rect -18 1000 18 1031
rect -18 -1031 18 -1000
rect -33 -1047 33 -1031
rect -33 -1081 -17 -1047
rect 17 -1081 33 -1047
rect -33 -1097 33 -1081
<< polycont >>
rect -17 1047 17 1081
rect -17 -1081 17 -1047
<< locali >>
rect -178 1149 -82 1183
rect 82 1149 178 1183
rect -178 1087 -144 1149
rect 144 1087 178 1149
rect -47 1047 -17 1081
rect 17 1047 47 1081
rect -64 988 -30 1004
rect -64 -1004 -30 -988
rect 30 988 64 1004
rect 30 -1004 64 -988
rect -47 -1081 -17 -1047
rect 17 -1081 47 -1047
rect -178 -1149 -144 -1087
rect 144 -1149 178 -1087
rect -178 -1183 -82 -1149
rect 82 -1183 178 -1149
<< viali >>
rect -17 1047 17 1081
rect -64 -988 -30 988
rect 30 -988 64 988
rect -17 -1081 17 -1047
<< metal1 >>
rect -29 1081 29 1087
rect -47 1047 -17 1081
rect 17 1047 47 1081
rect -29 1041 29 1047
rect -70 988 -24 1000
rect -70 -988 -64 988
rect -30 -988 -24 988
rect -70 -1000 -24 -988
rect 24 988 70 1000
rect 24 -988 30 988
rect 64 -988 70 988
rect 24 -1000 70 -988
rect -29 -1047 29 -1041
rect -47 -1081 -17 -1047
rect 17 -1081 47 -1047
rect -29 -1087 29 -1081
<< labels >>
rlabel nsubdiffcont 0 -1166 0 -1166 0 B
port 1 nsew
rlabel pdiffc -47 0 -47 0 0 D
port 2 nsew
rlabel pdiffc 47 0 47 0 0 S
port 3 nsew
rlabel polycont 0 1064 0 1064 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -161 -1166 161 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
