magic
tech sky130A
magscale 1 2
timestamp 1764202196
<< nwell >>
rect -246 -2555 246 2555
<< pmos >>
rect -50 936 50 2336
rect -50 -700 50 700
rect -50 -2336 50 -936
<< pdiff >>
rect -108 2324 -50 2336
rect -108 948 -96 2324
rect -62 948 -50 2324
rect -108 936 -50 948
rect 50 2324 108 2336
rect 50 948 62 2324
rect 96 948 108 2324
rect 50 936 108 948
rect -108 688 -50 700
rect -108 -688 -96 688
rect -62 -688 -50 688
rect -108 -700 -50 -688
rect 50 688 108 700
rect 50 -688 62 688
rect 96 -688 108 688
rect 50 -700 108 -688
rect -108 -948 -50 -936
rect -108 -2324 -96 -948
rect -62 -2324 -50 -948
rect -108 -2336 -50 -2324
rect 50 -948 108 -936
rect 50 -2324 62 -948
rect 96 -2324 108 -948
rect 50 -2336 108 -2324
<< pdiffc >>
rect -96 948 -62 2324
rect 62 948 96 2324
rect -96 -688 -62 688
rect 62 -688 96 688
rect -96 -2324 -62 -948
rect 62 -2324 96 -948
<< nsubdiff >>
rect -210 2485 -114 2519
rect 114 2485 210 2519
rect -210 2423 -176 2485
rect 176 2423 210 2485
rect -210 -2485 -176 -2423
rect 176 -2485 210 -2423
rect -210 -2519 -114 -2485
rect 114 -2519 210 -2485
<< nsubdiffcont >>
rect -114 2485 114 2519
rect -210 -2423 -176 2423
rect 176 -2423 210 2423
rect -114 -2519 114 -2485
<< poly >>
rect -50 2417 50 2433
rect -50 2383 -34 2417
rect 34 2383 50 2417
rect -50 2336 50 2383
rect -50 889 50 936
rect -50 855 -34 889
rect 34 855 50 889
rect -50 839 50 855
rect -50 781 50 797
rect -50 747 -34 781
rect 34 747 50 781
rect -50 700 50 747
rect -50 -747 50 -700
rect -50 -781 -34 -747
rect 34 -781 50 -747
rect -50 -797 50 -781
rect -50 -855 50 -839
rect -50 -889 -34 -855
rect 34 -889 50 -855
rect -50 -936 50 -889
rect -50 -2383 50 -2336
rect -50 -2417 -34 -2383
rect 34 -2417 50 -2383
rect -50 -2433 50 -2417
<< polycont >>
rect -34 2383 34 2417
rect -34 855 34 889
rect -34 747 34 781
rect -34 -781 34 -747
rect -34 -889 34 -855
rect -34 -2417 34 -2383
<< locali >>
rect -210 2485 -114 2519
rect 114 2485 210 2519
rect -210 2423 -176 2485
rect 176 2423 210 2485
rect -50 2383 -34 2417
rect 34 2383 50 2417
rect -96 2324 -62 2340
rect -96 932 -62 948
rect 62 2324 96 2340
rect 62 932 96 948
rect -50 855 -34 889
rect 34 855 50 889
rect -50 747 -34 781
rect 34 747 50 781
rect -96 688 -62 704
rect -96 -704 -62 -688
rect 62 688 96 704
rect 62 -704 96 -688
rect -50 -781 -34 -747
rect 34 -781 50 -747
rect -50 -889 -34 -855
rect 34 -889 50 -855
rect -96 -948 -62 -932
rect -96 -2340 -62 -2324
rect 62 -948 96 -932
rect 62 -2340 96 -2324
rect -50 -2417 -34 -2383
rect 34 -2417 50 -2383
rect -210 -2485 -176 -2423
rect 176 -2485 210 -2423
rect -210 -2519 -114 -2485
rect 114 -2519 210 -2485
<< viali >>
rect -34 2383 34 2417
rect -96 948 -62 2324
rect 62 948 96 2324
rect -34 855 34 889
rect -34 747 34 781
rect -96 -688 -62 688
rect 62 -688 96 688
rect -34 -781 34 -747
rect -34 -889 34 -855
rect -96 -2324 -62 -948
rect 62 -2324 96 -948
rect -34 -2417 34 -2383
<< metal1 >>
rect -46 2417 46 2423
rect -46 2383 -34 2417
rect 34 2383 46 2417
rect -46 2377 46 2383
rect -102 2324 -56 2336
rect -102 948 -96 2324
rect -62 948 -56 2324
rect -102 936 -56 948
rect 56 2324 102 2336
rect 56 948 62 2324
rect 96 948 102 2324
rect 56 936 102 948
rect -46 889 46 895
rect -46 855 -34 889
rect 34 855 46 889
rect -46 849 46 855
rect -46 781 46 787
rect -46 747 -34 781
rect 34 747 46 781
rect -46 741 46 747
rect -102 688 -56 700
rect -102 -688 -96 688
rect -62 -688 -56 688
rect -102 -700 -56 -688
rect 56 688 102 700
rect 56 -688 62 688
rect 96 -688 102 688
rect 56 -700 102 -688
rect -46 -747 46 -741
rect -46 -781 -34 -747
rect 34 -781 46 -747
rect -46 -787 46 -781
rect -46 -855 46 -849
rect -46 -889 -34 -855
rect 34 -889 46 -855
rect -46 -895 46 -889
rect -102 -948 -56 -936
rect -102 -2324 -96 -948
rect -62 -2324 -56 -948
rect -102 -2336 -56 -2324
rect 56 -948 102 -936
rect 56 -2324 62 -948
rect 96 -2324 102 -948
rect 56 -2336 102 -2324
rect -46 -2383 46 -2377
rect -46 -2417 -34 -2383
rect 34 -2417 46 -2383
rect -46 -2423 46 -2417
<< labels >>
rlabel nsubdiffcont 0 -2502 0 -2502 0 B
port 31 nsew
rlabel pdiffc -79 -1636 -79 -1636 0 D0
port 32 nsew
rlabel pdiffc 79 -1636 79 -1636 0 S0
port 33 nsew
rlabel polycont 0 -872 0 -872 0 G0
port 34 nsew
rlabel pdiffc -79 0 -79 0 0 D1
port 35 nsew
rlabel pdiffc 79 0 79 0 0 S1
port 36 nsew
rlabel polycont 0 764 0 764 0 G1
port 37 nsew
rlabel pdiffc -79 1636 -79 1636 0 D2
port 38 nsew
rlabel pdiffc 79 1636 79 1636 0 S2
port 39 nsew
rlabel polycont 0 2400 0 2400 0 G2
port 40 nsew
<< properties >>
string FIXED_BBOX -193 -2502 193 2502
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7 l 0.5 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
