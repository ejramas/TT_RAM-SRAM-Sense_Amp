magic
tech sky130A
magscale 1 2
timestamp 1764449767
<< nwell >>
rect -404 -919 404 919
<< pmos >>
rect -208 -700 -108 700
rect -50 -700 50 700
rect 108 -700 208 700
<< pdiff >>
rect -266 688 -208 700
rect -266 -688 -254 688
rect -220 -688 -208 688
rect -266 -700 -208 -688
rect -108 688 -50 700
rect -108 -688 -96 688
rect -62 -688 -50 688
rect -108 -700 -50 -688
rect 50 688 108 700
rect 50 -688 62 688
rect 96 -688 108 688
rect 50 -700 108 -688
rect 208 688 266 700
rect 208 -688 220 688
rect 254 -688 266 688
rect 208 -700 266 -688
<< pdiffc >>
rect -254 -688 -220 688
rect -96 -688 -62 688
rect 62 -688 96 688
rect 220 -688 254 688
<< nsubdiff >>
rect -368 849 -272 883
rect 272 849 368 883
rect -368 787 -334 849
rect 334 787 368 849
rect -368 -849 -334 -787
rect 334 -849 368 -787
rect -368 -883 -272 -849
rect 272 -883 368 -849
<< nsubdiffcont >>
rect -272 849 272 883
rect -368 -787 -334 787
rect 334 -787 368 787
rect -272 -883 272 -849
<< poly >>
rect -208 781 -108 797
rect -208 747 -192 781
rect -124 747 -108 781
rect -208 700 -108 747
rect -50 781 50 797
rect -50 747 -34 781
rect 34 747 50 781
rect -50 700 50 747
rect 108 781 208 797
rect 108 747 124 781
rect 192 747 208 781
rect 108 700 208 747
rect -208 -747 -108 -700
rect -208 -781 -192 -747
rect -124 -781 -108 -747
rect -208 -797 -108 -781
rect -50 -747 50 -700
rect -50 -781 -34 -747
rect 34 -781 50 -747
rect -50 -797 50 -781
rect 108 -747 208 -700
rect 108 -781 124 -747
rect 192 -781 208 -747
rect 108 -797 208 -781
<< polycont >>
rect -192 747 -124 781
rect -34 747 34 781
rect 124 747 192 781
rect -192 -781 -124 -747
rect -34 -781 34 -747
rect 124 -781 192 -747
<< locali >>
rect -368 849 -272 883
rect 272 849 368 883
rect -368 787 -334 849
rect 334 787 368 849
rect -237 747 -192 781
rect -124 747 -34 781
rect 34 747 124 781
rect 192 747 237 781
rect -254 688 -220 704
rect -254 -704 -220 -688
rect -96 688 -62 704
rect -96 -704 -62 -688
rect 62 688 96 704
rect 62 -704 96 -688
rect 220 688 254 704
rect 220 -704 254 -688
rect -237 -781 -192 -747
rect -124 -781 -34 -747
rect 34 -781 124 -747
rect 192 -781 237 -747
rect -368 -849 -334 -787
rect 334 -849 368 -787
rect -368 -883 -272 -849
rect 272 -883 368 -849
<< viali >>
rect -192 747 -124 781
rect -34 747 34 781
rect 124 747 192 781
rect -254 -688 -220 688
rect -96 -688 -62 688
rect 62 -688 96 688
rect 220 -688 254 688
rect -192 -781 -124 -747
rect -34 -781 34 -747
rect 124 -781 192 -747
<< metal1 >>
rect -204 781 -112 787
rect -46 781 46 787
rect 112 781 204 787
rect -237 747 -192 781
rect -124 747 -34 781
rect 34 747 124 781
rect 192 747 237 781
rect -204 741 -112 747
rect -46 741 46 747
rect 112 741 204 747
rect -260 688 -214 700
rect -260 -688 -254 688
rect -220 -688 -214 688
rect -260 -700 -214 -688
rect -102 688 -56 700
rect -102 -688 -96 688
rect -62 -688 -56 688
rect -102 -700 -56 -688
rect 56 688 102 700
rect 56 -688 62 688
rect 96 -688 102 688
rect 56 -700 102 -688
rect 214 688 260 700
rect 214 -688 220 688
rect 254 -688 260 688
rect 214 -700 260 -688
rect -204 -747 -112 -741
rect -46 -747 46 -741
rect 112 -747 204 -741
rect -237 -781 -192 -747
rect -124 -781 -34 -747
rect 34 -781 124 -747
rect 192 -781 237 -747
rect -204 -787 -112 -781
rect -46 -787 46 -781
rect 112 -787 204 -781
<< labels >>
rlabel nsubdiffcont 0 -866 0 -866 0 B
port 1 nsew
rlabel pdiffc -237 0 -237 0 0 D0
port 2 nsew
rlabel polycont -158 764 -158 764 0 G
port 3 nsew
rlabel pdiffc -79 0 -79 0 0 S1
port 4 nsew
rlabel polycont 0 764 0 764 0 G
port 3 nsew
rlabel pdiffc 79 0 79 0 0 D2
port 5 nsew
rlabel pdiffc 237 0 237 0 0 S2
port 6 nsew
rlabel polycont 158 764 158 764 0 G
port 3 nsew
<< properties >>
string FIXED_BBOX -351 -866 351 866
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7 l 0.5 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
