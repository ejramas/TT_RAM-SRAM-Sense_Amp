magic
tech sky130A
magscale 1 2
timestamp 1764202196
<< error_p >>
rect -29 590 29 596
rect -29 556 -17 590
rect -29 550 29 556
rect -29 280 29 286
rect -29 246 -17 280
rect -29 240 29 246
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect -29 -178 29 -172
rect -29 -246 29 -240
rect -29 -280 -17 -246
rect -29 -286 29 -280
rect -29 -556 29 -550
rect -29 -590 -17 -556
rect -29 -596 29 -590
<< pwell >>
rect -214 -728 214 728
<< nmos >>
rect -18 318 18 518
rect -18 -100 18 100
rect -18 -518 18 -318
<< ndiff >>
rect -76 506 -18 518
rect -76 330 -64 506
rect -30 330 -18 506
rect -76 318 -18 330
rect 18 506 76 518
rect 18 330 30 506
rect 64 330 76 506
rect 18 318 76 330
rect -76 88 -18 100
rect -76 -88 -64 88
rect -30 -88 -18 88
rect -76 -100 -18 -88
rect 18 88 76 100
rect 18 -88 30 88
rect 64 -88 76 88
rect 18 -100 76 -88
rect -76 -330 -18 -318
rect -76 -506 -64 -330
rect -30 -506 -18 -330
rect -76 -518 -18 -506
rect 18 -330 76 -318
rect 18 -506 30 -330
rect 64 -506 76 -330
rect 18 -518 76 -506
<< ndiffc >>
rect -64 330 -30 506
rect 30 330 64 506
rect -64 -88 -30 88
rect 30 -88 64 88
rect -64 -506 -30 -330
rect 30 -506 64 -330
<< psubdiff >>
rect -178 658 -82 692
rect 82 658 178 692
rect -178 596 -144 658
rect 144 596 178 658
rect -178 -658 -144 -596
rect 144 -658 178 -596
rect -178 -692 -82 -658
rect 82 -692 178 -658
<< psubdiffcont >>
rect -82 658 82 692
rect -178 -596 -144 596
rect 144 -596 178 596
rect -82 -692 82 -658
<< poly >>
rect -33 590 33 606
rect -33 556 -17 590
rect 17 556 33 590
rect -33 540 33 556
rect -18 518 18 540
rect -18 296 18 318
rect -33 280 33 296
rect -33 246 -17 280
rect 17 246 33 280
rect -33 230 33 246
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -18 100 18 122
rect -18 -122 18 -100
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
rect -33 -246 33 -230
rect -33 -280 -17 -246
rect 17 -280 33 -246
rect -33 -296 33 -280
rect -18 -318 18 -296
rect -18 -540 18 -518
rect -33 -556 33 -540
rect -33 -590 -17 -556
rect 17 -590 33 -556
rect -33 -606 33 -590
<< polycont >>
rect -17 556 17 590
rect -17 246 17 280
rect -17 138 17 172
rect -17 -172 17 -138
rect -17 -280 17 -246
rect -17 -590 17 -556
<< locali >>
rect -178 658 -82 692
rect 82 658 178 692
rect -178 596 -144 658
rect 144 596 178 658
rect -33 556 -17 590
rect 17 556 33 590
rect -64 506 -30 522
rect -64 314 -30 330
rect 30 506 64 522
rect 30 314 64 330
rect -33 246 -17 280
rect 17 246 33 280
rect -33 138 -17 172
rect 17 138 33 172
rect -64 88 -30 104
rect -64 -104 -30 -88
rect 30 88 64 104
rect 30 -104 64 -88
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -280 -17 -246
rect 17 -280 33 -246
rect -64 -330 -30 -314
rect -64 -522 -30 -506
rect 30 -330 64 -314
rect 30 -522 64 -506
rect -33 -590 -17 -556
rect 17 -590 33 -556
rect -178 -658 -144 -596
rect 144 -658 178 -596
rect -178 -692 -82 -658
rect 82 -692 178 -658
<< viali >>
rect -17 556 17 590
rect -64 330 -30 506
rect 30 330 64 506
rect -17 246 17 280
rect -17 138 17 172
rect -64 -88 -30 88
rect 30 -88 64 88
rect -17 -172 17 -138
rect -17 -280 17 -246
rect -64 -506 -30 -330
rect 30 -506 64 -330
rect -17 -590 17 -556
<< metal1 >>
rect -29 590 29 596
rect -29 556 -17 590
rect 17 556 29 590
rect -29 550 29 556
rect -70 506 -24 518
rect -70 330 -64 506
rect -30 330 -24 506
rect -70 318 -24 330
rect 24 506 70 518
rect 24 330 30 506
rect 64 330 70 506
rect 24 318 70 330
rect -29 280 29 286
rect -29 246 -17 280
rect 17 246 29 280
rect -29 240 29 246
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -70 88 -24 100
rect -70 -88 -64 88
rect -30 -88 -24 88
rect -70 -100 -24 -88
rect 24 88 70 100
rect 24 -88 30 88
rect 64 -88 70 88
rect 24 -100 70 -88
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
rect -29 -246 29 -240
rect -29 -280 -17 -246
rect 17 -280 29 -246
rect -29 -286 29 -280
rect -70 -330 -24 -318
rect -70 -506 -64 -330
rect -30 -506 -24 -330
rect -70 -518 -24 -506
rect 24 -330 70 -318
rect 24 -506 30 -330
rect 64 -506 70 -330
rect 24 -518 70 -506
rect -29 -556 29 -550
rect -29 -590 -17 -556
rect 17 -590 29 -556
rect -29 -596 29 -590
<< labels >>
rlabel psubdiffcont 0 -675 0 -675 0 B
port 1 nsew
rlabel ndiffc -47 -418 -47 -418 0 D0
port 2 nsew
rlabel ndiffc 47 -418 47 -418 0 S0
port 3 nsew
rlabel polycont 0 -263 0 -263 0 G0
port 4 nsew
rlabel ndiffc -47 0 -47 0 0 D1
port 5 nsew
rlabel ndiffc 47 0 47 0 0 S1
port 6 nsew
rlabel polycont 0 155 0 155 0 G1
port 7 nsew
rlabel ndiffc -47 418 -47 418 0 D2
port 8 nsew
rlabel ndiffc 47 418 47 418 0 S2
port 9 nsew
rlabel polycont 0 573 0 573 0 G2
port 10 nsew
<< properties >>
string FIXED_BBOX -161 -675 161 675
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.18 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
