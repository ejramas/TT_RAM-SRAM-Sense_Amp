magic
tech sky130A
magscale 1 2
timestamp 1764871086
<< viali >>
rect 1940 6180 2000 6280
rect 4140 6220 4220 6320
rect 1060 5940 1160 6040
rect 4820 5880 4900 5960
rect 1520 5480 1580 5540
rect 4380 5420 4440 5480
rect 4120 4760 4180 4820
rect 1520 4600 1580 4660
rect 3620 4560 3680 4620
rect 2680 4240 2740 4300
rect 3380 4240 3440 4300
rect 2680 3720 2740 3780
rect 3320 3720 3380 3780
<< metal1 >>
rect 4960 7360 5100 7380
rect 860 7320 1020 7340
rect 860 7200 880 7320
rect 1000 7200 1020 7320
rect 860 7120 1020 7200
rect 4960 7280 4980 7360
rect 5080 7280 5100 7360
rect 4960 7180 5100 7280
rect 5000 6760 5020 6800
rect 960 6600 2560 6720
rect 3580 6620 5020 6760
rect 5080 6620 5120 6760
rect 1580 6440 1780 6460
rect 1820 6440 1940 6600
rect 1580 6340 1600 6440
rect 1680 6340 1780 6440
rect 1580 6320 1780 6340
rect 1920 6280 2020 6360
rect 2060 6340 2120 6460
rect 4020 6380 4080 6500
rect 4200 6460 4320 6620
rect 4360 6480 4540 6500
rect 4360 6400 4440 6480
rect 4520 6400 4540 6480
rect 4960 6440 5020 6480
rect 5080 6440 5100 6480
rect 1920 6180 1940 6280
rect 2000 6180 2020 6280
rect 700 6040 920 6060
rect 700 5940 720 6040
rect 800 5940 920 6040
rect 700 5920 920 5940
rect 1040 6040 1180 6060
rect 1040 5940 1060 6040
rect 1160 5940 1180 6040
rect 1040 5920 1180 5940
rect 860 2980 1020 3060
rect 860 2880 880 2980
rect 1000 2880 1020 2980
rect 1260 3020 1340 6100
rect 1920 6060 2020 6180
rect 4120 6320 4240 6400
rect 4360 6380 4540 6400
rect 4120 6220 4140 6320
rect 4220 6220 4240 6320
rect 4120 6060 4240 6220
rect 1920 5940 4240 6060
rect 1500 5880 4240 5940
rect 1500 5840 4460 5880
rect 1500 5540 1600 5840
rect 1920 5780 4460 5840
rect 1920 5720 4240 5780
rect 1920 5660 1940 5720
rect 2020 5660 2520 5720
rect 2600 5660 3540 5720
rect 3620 5660 4120 5720
rect 4200 5660 4240 5720
rect 1920 5640 4240 5660
rect 1720 5540 1940 5600
rect 2020 5540 2060 5600
rect 1500 5480 1520 5540
rect 1580 5480 1600 5540
rect 1500 5460 1600 5480
rect 1720 5440 1740 5500
rect 1820 5440 2060 5500
rect 1720 5340 1940 5400
rect 2020 5340 2060 5400
rect 1720 5220 1740 5280
rect 1820 5220 2060 5280
rect 2100 5260 2240 5560
rect 2300 5540 2520 5600
rect 2600 5540 2620 5600
rect 2300 5440 2320 5500
rect 2400 5440 2620 5500
rect 2300 5340 2520 5400
rect 2600 5340 2620 5400
rect 2300 5240 2320 5300
rect 2400 5240 2620 5300
rect 2660 5260 3300 5560
rect 3340 5540 3540 5600
rect 3620 5540 3660 5600
rect 3340 5440 3360 5500
rect 3440 5440 3660 5500
rect 3340 5340 3540 5400
rect 3620 5340 3660 5400
rect 2660 5180 2820 5260
rect 3340 5240 3360 5300
rect 3440 5240 3660 5300
rect 3720 5260 3860 5560
rect 3920 5540 4120 5600
rect 4200 5540 4240 5600
rect 3920 5440 3940 5500
rect 4020 5440 4240 5500
rect 4360 5480 4460 5780
rect 4360 5420 4380 5480
rect 4440 5420 4460 5480
rect 4360 5400 4460 5420
rect 3920 5340 4120 5400
rect 4200 5340 4240 5400
rect 3920 5240 3940 5300
rect 4020 5240 4240 5300
rect 1720 5160 2820 5180
rect 1720 5100 1740 5160
rect 1820 5100 2320 5160
rect 2400 5100 2820 5160
rect 1720 5020 2820 5100
rect 1480 4920 1740 4940
rect 1480 4860 1640 4920
rect 1720 4860 1740 4920
rect 1480 4840 1740 4860
rect 1480 4660 1600 4840
rect 1480 4600 1520 4660
rect 1580 4600 1600 4660
rect 1480 4580 1600 4600
rect 1480 4480 1680 4580
rect 1920 4560 2040 4580
rect 2660 4560 2820 5020
rect 3340 4920 4560 4940
rect 3340 4860 3360 4920
rect 3440 4860 4560 4920
rect 3340 4840 4560 4860
rect 4100 4820 4200 4840
rect 4100 4760 4120 4820
rect 4180 4760 4200 4820
rect 4100 4740 4200 4760
rect 3240 4620 3360 4640
rect 3240 4560 3260 4620
rect 3340 4560 3360 4620
rect 3600 4620 3700 4640
rect 3600 4560 3620 4620
rect 3680 4560 3700 4620
rect 4440 4560 4560 4840
rect 1920 4500 1940 4560
rect 2020 4500 2040 4560
rect 3240 4540 3440 4560
rect 3600 4540 3700 4560
rect 4000 4540 4120 4560
rect 1920 4480 2040 4500
rect 3380 4440 3440 4540
rect 4000 4480 4020 4540
rect 4100 4480 4120 4540
rect 4000 4460 4120 4480
rect 4360 4540 4560 4560
rect 4360 4480 4460 4540
rect 4540 4480 4560 4540
rect 4360 4460 4560 4480
rect 2680 4360 3440 4440
rect 2680 4320 2740 4360
rect 3380 4320 3440 4360
rect 2660 4300 2760 4320
rect 2660 4240 2680 4300
rect 2740 4240 2760 4300
rect 2660 4220 2760 4240
rect 3360 4300 3460 4320
rect 3360 4240 3380 4300
rect 3440 4240 3460 4300
rect 3360 4220 3460 4240
rect 2680 4180 2740 4220
rect 3380 4180 3440 4220
rect 2340 4100 2560 4140
rect 3500 4100 3640 4140
rect 2340 3640 2380 4100
rect 2660 3860 2760 4060
rect 3300 3860 3400 4060
rect 2660 3840 2900 3860
rect 2660 3780 2800 3840
rect 2880 3780 2900 3840
rect 2660 3720 2680 3780
rect 2740 3760 2900 3780
rect 3160 3840 3400 3860
rect 3160 3780 3180 3840
rect 3260 3780 3400 3840
rect 3160 3760 3320 3780
rect 2740 3720 2760 3760
rect 2660 3660 2760 3720
rect 3300 3720 3320 3760
rect 3380 3720 3400 3780
rect 3300 3660 3400 3720
rect 2160 3560 2380 3640
rect 1760 3520 1880 3540
rect 1760 3460 1780 3520
rect 1860 3460 1880 3520
rect 1760 3440 1880 3460
rect 2260 3520 2380 3560
rect 3600 3640 3640 4100
rect 3600 3560 3900 3640
rect 2260 3460 2280 3520
rect 2360 3460 2380 3520
rect 1940 3020 1980 3140
rect 2260 3120 2380 3460
rect 2640 3520 2760 3540
rect 2640 3460 2660 3520
rect 2740 3460 2760 3520
rect 2640 3440 2760 3460
rect 3280 3520 3400 3540
rect 3280 3460 3300 3520
rect 3380 3460 3400 3520
rect 3280 3440 3400 3460
rect 3600 3520 3720 3560
rect 3600 3460 3620 3520
rect 3700 3460 3720 3520
rect 2640 3360 2760 3380
rect 2640 3300 2660 3360
rect 2740 3300 2760 3360
rect 2640 3280 2760 3300
rect 3300 3360 3420 3380
rect 3300 3300 3320 3360
rect 3400 3300 3420 3360
rect 3300 3280 3420 3300
rect 2260 3060 2280 3120
rect 2360 3080 2380 3120
rect 2640 3080 2780 3160
rect 2360 3060 2780 3080
rect 2260 3040 2780 3060
rect 1260 2960 1980 3020
rect 2840 2960 2880 3200
rect 1260 2920 2880 2960
rect 3180 2960 3220 3200
rect 3280 3060 3420 3160
rect 3600 3100 3720 3460
rect 4160 3520 4280 3540
rect 4160 3460 4180 3520
rect 4260 3460 4280 3520
rect 4160 3440 4280 3460
rect 3600 3060 3620 3100
rect 3280 3040 3620 3060
rect 3700 3040 3720 3100
rect 3280 3020 3720 3040
rect 4060 3020 4100 3140
rect 4620 3020 4700 6120
rect 4800 5960 4920 5980
rect 4800 5880 4820 5960
rect 4900 5880 4920 5960
rect 4800 5860 4920 5880
rect 5040 5960 5160 5980
rect 5040 5880 5060 5960
rect 5140 5880 5160 5960
rect 5040 5860 5160 5880
rect 4060 2960 4700 3020
rect 3180 2920 4700 2960
rect 4980 2960 5100 3120
rect 860 2860 1020 2880
rect 4980 2880 5000 2960
rect 5080 2880 5100 2960
rect 4980 2860 5100 2880
<< via1 >>
rect 880 7200 1000 7320
rect 4980 7280 5080 7360
rect 1600 6340 1680 6440
rect 4440 6400 4520 6480
rect 720 5940 800 6040
rect 1060 5940 1160 6040
rect 880 2880 1000 2980
rect 1940 5660 2020 5720
rect 2520 5660 2600 5720
rect 3540 5660 3620 5720
rect 4120 5660 4200 5720
rect 1940 5540 2020 5600
rect 1740 5440 1820 5500
rect 1940 5340 2020 5400
rect 1740 5220 1820 5280
rect 2520 5540 2600 5600
rect 2320 5440 2400 5500
rect 2520 5340 2600 5400
rect 2320 5240 2400 5300
rect 3540 5540 3620 5600
rect 3360 5440 3440 5500
rect 3540 5340 3620 5400
rect 3360 5240 3440 5300
rect 4120 5540 4200 5600
rect 3940 5440 4020 5500
rect 4120 5340 4200 5400
rect 3940 5240 4020 5300
rect 1740 5100 1820 5160
rect 2320 5100 2400 5160
rect 1640 4860 1720 4920
rect 3360 4860 3440 4920
rect 3260 4560 3340 4620
rect 3620 4560 3680 4620
rect 1940 4500 2020 4560
rect 4020 4480 4100 4540
rect 4460 4480 4540 4540
rect 2800 3780 2880 3840
rect 3180 3780 3260 3840
rect 1780 3460 1860 3520
rect 2280 3460 2360 3520
rect 2660 3460 2740 3520
rect 3300 3460 3380 3520
rect 3620 3460 3700 3520
rect 2660 3300 2740 3360
rect 3320 3300 3400 3360
rect 2280 3060 2360 3120
rect 4180 3460 4260 3520
rect 3620 3040 3700 3100
rect 4840 5880 4900 5960
rect 5060 5880 5140 5960
rect 5000 2880 5080 2960
<< metal2 >>
rect 4420 7360 5100 7380
rect 860 7320 1700 7340
rect 860 7200 880 7320
rect 1000 7200 1700 7320
rect 860 7180 1700 7200
rect 1580 6440 1700 7180
rect 1580 6340 1600 6440
rect 1680 6340 1700 6440
rect 4420 7280 4980 7360
rect 5080 7280 5100 7360
rect 4420 7260 5100 7280
rect 4420 6480 4540 7260
rect 4420 6400 4440 6480
rect 4520 6400 4540 6480
rect 4420 6380 4540 6400
rect 1580 6320 1700 6340
rect 700 6040 1260 6060
rect 700 5940 720 6040
rect 800 5940 1060 6040
rect 1160 6000 1260 6040
rect 1340 6020 4580 6060
rect 1340 6000 2900 6020
rect 1160 5940 2900 6000
rect 700 5920 2900 5940
rect 2980 5980 4580 6020
rect 2980 5960 5160 5980
rect 2980 5920 4840 5960
rect 4460 5880 4840 5920
rect 4900 5880 5060 5960
rect 5140 5880 5160 5960
rect 4460 5860 5160 5880
rect 1920 5720 2040 5740
rect 1920 5660 1940 5720
rect 2020 5660 2040 5720
rect 1920 5600 2040 5660
rect 1920 5540 1940 5600
rect 2020 5540 2040 5600
rect 1720 5500 1840 5520
rect 1720 5440 1740 5500
rect 1820 5440 1840 5500
rect 1720 5280 1840 5440
rect 1920 5400 2040 5540
rect 2500 5720 2620 5740
rect 2500 5660 2520 5720
rect 2600 5660 2620 5720
rect 2500 5600 2620 5660
rect 2500 5540 2520 5600
rect 2600 5540 2620 5600
rect 1920 5340 1940 5400
rect 2020 5340 2040 5400
rect 1920 5320 2040 5340
rect 2300 5500 2420 5520
rect 2300 5440 2320 5500
rect 2400 5440 2420 5500
rect 1720 5220 1740 5280
rect 1820 5220 1840 5280
rect 1720 5160 1840 5220
rect 1720 5100 1740 5160
rect 1820 5100 1840 5160
rect 1720 5080 1840 5100
rect 2300 5300 2420 5440
rect 2500 5400 2620 5540
rect 3520 5720 3640 5740
rect 3520 5660 3540 5720
rect 3620 5660 3640 5720
rect 3520 5600 3640 5660
rect 3520 5540 3540 5600
rect 3620 5540 3640 5600
rect 2500 5340 2520 5400
rect 2600 5340 2620 5400
rect 2500 5320 2620 5340
rect 3340 5500 3460 5520
rect 3340 5440 3360 5500
rect 3440 5440 3460 5500
rect 2300 5240 2320 5300
rect 2400 5240 2420 5300
rect 2300 5160 2420 5240
rect 2300 5100 2320 5160
rect 2400 5100 2420 5160
rect 2300 5080 2420 5100
rect 3340 5300 3460 5440
rect 3520 5400 3640 5540
rect 4100 5720 4220 5740
rect 4100 5660 4120 5720
rect 4200 5660 4220 5720
rect 4100 5600 4220 5660
rect 4100 5540 4120 5600
rect 4200 5540 4220 5600
rect 3520 5340 3540 5400
rect 3620 5340 3640 5400
rect 3520 5320 3640 5340
rect 3920 5500 4040 5520
rect 3920 5440 3940 5500
rect 4020 5440 4040 5500
rect 3340 5240 3360 5300
rect 3440 5240 3460 5300
rect 3340 5200 3460 5240
rect 3920 5300 4040 5440
rect 4100 5400 4220 5540
rect 4100 5340 4120 5400
rect 4200 5340 4220 5400
rect 4100 5320 4220 5340
rect 3920 5240 3940 5300
rect 4020 5240 4040 5300
rect 3920 5200 4040 5240
rect 3340 5120 4040 5200
rect 3340 4940 3460 5120
rect 1620 4920 3460 4940
rect 1620 4860 1640 4920
rect 1720 4860 3360 4920
rect 3440 4860 3460 4920
rect 4460 4860 4580 5860
rect 1620 4840 3460 4860
rect 1920 4560 2040 4840
rect 3660 4720 4580 4860
rect 3660 4660 3780 4720
rect 1920 4500 1940 4560
rect 2020 4500 2040 4560
rect 3240 4620 3780 4660
rect 3240 4560 3260 4620
rect 3340 4560 3620 4620
rect 3680 4560 3780 4620
rect 3240 4520 3780 4560
rect 4000 4540 4560 4560
rect 1920 4480 2040 4500
rect 4000 4480 4020 4540
rect 4100 4480 4460 4540
rect 4540 4480 4560 4540
rect 4000 4460 4560 4480
rect 2780 3840 2900 3860
rect 2780 3780 2800 3840
rect 2880 3780 2900 3840
rect 2780 3760 2900 3780
rect 2840 3740 2900 3760
rect 3160 3840 3280 3860
rect 3160 3780 3180 3840
rect 3260 3780 3280 3840
rect 3160 3760 3280 3780
rect 3160 3740 3220 3760
rect 2840 3680 3220 3740
rect 1760 3520 2760 3540
rect 1760 3460 1780 3520
rect 1860 3460 2280 3520
rect 2360 3460 2660 3520
rect 2740 3460 2760 3520
rect 1760 3440 2760 3460
rect 2840 3380 2900 3680
rect 2640 3360 2900 3380
rect 2640 3300 2660 3360
rect 2740 3300 2900 3360
rect 2640 3280 2900 3300
rect 3160 3380 3220 3680
rect 3280 3520 4280 3540
rect 3280 3460 3300 3520
rect 3380 3460 3620 3520
rect 3700 3460 4180 3520
rect 4260 3460 4280 3520
rect 3280 3440 4280 3460
rect 3160 3360 3420 3380
rect 3160 3300 3320 3360
rect 3400 3300 3420 3360
rect 3160 3280 3420 3300
rect 2260 3120 2380 3140
rect 2260 3060 2280 3120
rect 2360 3060 2380 3120
rect 2260 3000 2380 3060
rect 860 2980 2380 3000
rect 860 2880 880 2980
rect 1000 2880 2380 2980
rect 860 2860 2380 2880
rect 3600 3100 3720 3120
rect 3600 3040 3620 3100
rect 3700 3040 3720 3100
rect 3600 2980 3720 3040
rect 3600 2960 5100 2980
rect 3600 2880 5000 2960
rect 5080 2880 5100 2960
rect 3600 2860 5100 2880
use sky130_fd_pr__nfet_01v8_2BLVHV  sky130_fd_pr__nfet_01v8_2BLVHV_0
timestamp 1764449767
transform 0 1 2710 -1 0 4114
box -214 -310 214 310
use sky130_fd_pr__nfet_01v8_2BLVHV  sky130_fd_pr__nfet_01v8_2BLVHV_1
timestamp 1764449767
transform 0 1 3350 -1 0 4114
box -214 -310 214 310
use sky130_fd_pr__nfet_01v8_49EKDV  sky130_fd_pr__nfet_01v8_49EKDV_0
timestamp 1764737709
transform -1 0 938 0 -1 5090
box -218 -2210 218 2210
use sky130_fd_pr__nfet_01v8_49EKDV  sky130_fd_pr__nfet_01v8_49EKDV_1
timestamp 1764737709
transform -1 0 5038 0 -1 5150
box -218 -2210 218 2210
use sky130_fd_pr__nfet_01v8_K8VX6U  sky130_fd_pr__nfet_01v8_K8VX6U_0
timestamp 1764636235
transform 0 1 3350 -1 0 3404
box -404 -310 404 310
use sky130_fd_pr__nfet_01v8_K8VX6U  sky130_fd_pr__nfet_01v8_K8VX6U_1
timestamp 1764636235
transform 0 1 2710 -1 0 3404
box -404 -310 404 310
use sky130_fd_pr__pfet_01v8_L3H7YA  sky130_fd_pr__pfet_01v8_L3H7YA_0
timestamp 1764451811
transform 0 1 3791 -1 0 5411
box -311 -671 311 671
use sky130_fd_pr__pfet_01v8_L3H7YA  sky130_fd_pr__pfet_01v8_L3H7YA_1
timestamp 1764451811
transform 0 1 2171 -1 0 5411
box -311 -671 311 671
use sky130_fd_pr__pfet_01v8_TGVDXL  sky130_fd_pr__pfet_01v8_TGVDXL_0
timestamp 1764449767
transform 1 0 1904 0 1 3919
box -404 -919 404 919
use sky130_fd_pr__pfet_01v8_TGVDXL  sky130_fd_pr__pfet_01v8_TGVDXL_1
timestamp 1764449767
transform 1 0 4144 0 1 3919
box -404 -919 404 919
use sky130_fd_pr__pfet_01v8_VKLFMA  sky130_fd_pr__pfet_01v8_VKLFMA_0
timestamp 1764737709
transform 0 1 4219 -1 0 6438
box -218 -319 218 319
use sky130_fd_pr__pfet_01v8_VKLFMA  sky130_fd_pr__pfet_01v8_VKLFMA_1
timestamp 1764737709
transform 0 1 1919 -1 0 6398
box -218 -319 218 319
use sky130_fd_pr__res_xhigh_po_0p35_RJXVHX  sky130_fd_pr__res_xhigh_po_0p35_RJXVHX_0
timestamp 1764638150
transform 0 -1 3051 1 0 4581
box -201 -651 201 651
<< labels >>
rlabel metal2 4500 5940 4540 5980 1 GND
port 2 n
rlabel metal1 2920 5960 2960 6000 1 VDD
port 1 n
rlabel metal1 4640 6040 4680 6080 1 bitline_n
port 4 n
rlabel metal1 1280 6020 1320 6060 1 bitline_p
port 3 n
rlabel metal1 2940 5380 2980 5420 1 comgate
port 7 n
rlabel metal1 3540 4880 3580 4920 1 vdp
port 8 n
rlabel metal1 2700 3860 2720 3880 1 vsp
port 9 n
rlabel metal1 3620 6660 3660 6700 1 new_out_n
port 6 n
rlabel metal1 2500 6640 2540 6680 1 new_out_p
port 5 n
<< end >>
